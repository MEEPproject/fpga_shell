// Here is the RTL needed in the EA to set the PCIe AXI communication
