    input          qsfp1_ref_clk_n ,
    input          qsfp1_ref_clk_p ,
    input   [0:0]  qsfp1_1x_grx_n ,
    input   [0:0]  qsfp1_1x_grx_p ,
    output  [0:0]  qsfp1_1x_gtx_n ,
    output  [0:0]  qsfp1_1x_gtx_p ,
    output         qsfp1_oe_b ,
    output         qsfp1_fs ,

