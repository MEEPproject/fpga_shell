# Place here a message that gets included in the automatically top shell file
