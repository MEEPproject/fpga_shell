
axi4_awready   
axi4_awvalid   
axi4_awid      
axi4_awuser    
axi4_awaddr    
axi4_awprot    
axi4_awqos     
axi4_awregion  
axi4_awlen     
axi4_awsize    
axi4_awburst   
axi4_awlock    
axi4_awcache   

axi4_wready    
axi4_wvalid    
axi4_wdata     
axi4_wuser     
axi4_wstrb     
axi4_wlast     

axi4_bready    
axi4_bvalid    
axi4_bid       
axi4_buser     
axi4_bresp     

axi4_arready   
axi4_arvalid   
axi4_arid      
axi4_aruser    
axi4_araddr    
axi4_arprot    
axi4_arqos     
axi4_arregion  
axi4_arlen     
axi4_arsize    
axi4_arburst   
axi4_arlock    
axi4_arcache   

axi4_rready    
axi4_rvalid    
axi4_rid       
axi4_ruser     
axi4_rresp     
axi4_rdata     
axi4_rlast     

