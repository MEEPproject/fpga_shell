    // DDR4
    output [0:0]  ddr4_sdram_c0_act_n   ,
    output [16:0] ddr4_sdram_c0_adr     ,
    output [1:0]  ddr4_sdram_c0_ba      ,
    output [1:0]  ddr4_sdram_c0_bg      ,
    output [0:0]  ddr4_sdram_c0_ck_c    ,
    output [0:0]  ddr4_sdram_c0_ck_t    ,
    output [0:0]  ddr4_sdram_c0_cke     ,
    output [0:0]  ddr4_sdram_c0_cs_n    ,
    inout  [71:0] ddr4_sdram_c0_dq      ,
    inout  [17:0] ddr4_sdram_c0_dqs_c   ,
    inout  [17:0] ddr4_sdram_c0_dqs_t   ,
    output [0:0]  ddr4_sdram_c0_odt     ,
    output [0:0]  ddr4_sdram_c0_par     ,
    output [0:0]  ddr4_sdram_c0_reset_n ,
