
axilite_awready   
axilite_awvalid     
axilite_awaddr    

axilite_wready    
axilite_wvalid    
axilite_wdata        
axilite_wstrb     
   
axilite_bready    
axilite_bvalid       
axilite_bresp     

axilite_arready   
axilite_arvalid     
axilite_araddr    

axilite_rready    
axilite_rvalid        
axilite_rresp     
axilite_rdata     
 

