    // UART
    input         rs232_rxd  ,
    output        rs232_txd  ,
