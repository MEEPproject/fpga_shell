
axiL_awready   
axiL_awvalid     
axiL_awaddr    

axiL_wready    
axiL_wvalid    
axiL_wdata        
axiL_wstrb     
   
axiL_bready    
axiL_bvalid       
axiL_bresp     

axiL_arready   
axiL_arvalid     
axiL_araddr    

axiL_rready    
axiL_rvalid        
axiL_rresp     
axiL_rdata     
 

