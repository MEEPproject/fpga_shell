    input          qsfp_ref_clk_n ,
    input          qsfp_ref_clk_p ,
    input   [3:0]  qsfp_4x_grx_n ,
    input   [3:0]  qsfp_4x_grx_p ,
    output  [3:0]  qsfp_4x_gtx_n ,
    output  [3:0]  qsfp_4x_gtx_p ,
