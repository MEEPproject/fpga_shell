// This is an RTL template useful when the 10Gb Ethernet IP is used
