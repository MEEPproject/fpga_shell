    // PCI express
	input         pcie_refclk_clk_n    ,
    input         pcie_refclk_clk_p    ,
    input         pcie_perstn          ,		
    input  [15:0] pci_express_x16_rxn  ,
    input  [15:0] pci_express_x16_rxp  ,
    output [15:0] pci_express_x16_txn  ,
    output [15:0] pci_express_x16_txp  ,