    // Main input clock
    input         sysclk0_clk_n  ,
    input         sysclk0_clk_p  ,
    // Secondary clock
    input         sysclk1_clk_n  ,
    input         sysclk1_clk_p  , 
    // Secondary clock
    //input         sysclk3_clk_n  ,
    //input         sysclk3_clk_p  ,	
	// system reset - CPU_RESET L30
    input         resetn  ,
