    input          qsfp0_ref_clk_n ,
    input          qsfp0_ref_clk_p ,
    input   [0:0]  qsfp0_1x_grx_n ,
    input   [0:0]  qsfp0_1x_grx_p ,
    output  [0:0]  qsfp0_1x_gtx_n ,
    output  [0:0]  qsfp0_1x_gtx_p ,
    output         qsfp0_oe_b ,
    output         qsfp0_fs ,

